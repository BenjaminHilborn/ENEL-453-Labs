-- PIN NUMBERS
-- Clock: B8
-- Push button: G12 OR C11 OR M4 OR A7
-- Anodes: 
--	AN0: F12
--	AN1: J12
--	AN2: M13
--	AN3: K14
-- Cathodes: 
--	CA: L14
--	CB: H12
--	CC: N14
--	CD: N11
--	CE: P12
--	CF: L13
--	CG: M12
-- Decimal point: N13
-- Slide switch: P11 OR L3 OR K3 OR B4 OR G3 OR F3 OR E2 OR N3